module assembler_Op (
    // INPUT
    input wire [31:0] PC_out,
    input wire [4:0] RS, RT,

    //OUTPUT
    output wire [31:0] SH_out,
    output wire [31:0] SB_out,
    output wire [31:0] S_out,
);
    assign SH_out = /*      */
    assign SB_out = /*      */
    assign S_out = /*       */
endmodule