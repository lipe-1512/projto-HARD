module assembler_Op (
    input wire [31:0] PC_out,
);
    
endmodule